module verilog_module();





	initial begin 


	end




endmodule;