// this is  top level module that works to instantiate other modules
module verilog_module();


mod1 m1();
mod2 m2();


	




endmodule;

module mod1;

endmodule 


module mod2;


endmodule