`include "../8_D_flip_flop/D_FF.v"

module shift_reg(
	input clk, 
	input D,
	output k,
	input rstn);

	






endmodule