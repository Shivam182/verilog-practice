module mm;

initial begin 

$display("hello i am shivam");

end

endmodule
