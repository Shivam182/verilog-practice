module hello(M,N);

    input M;
    output N;

    assign N = M;



endmodule